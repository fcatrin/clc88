parameter VGA_MODE_640x480   = 2'b01;
parameter VGA_MODE_800x600   = 2'b10;
parameter VGA_MODE_1920x1080 = 2'b11;