parameter OP_NOP      = 0;
parameter OP_UPDATE   = 1;
parameter OP_AND      = 2;
parameter OP_OR       = 3;
parameter OP_EOR      = 4;
parameter OP_ADD      = 5;
parameter OP_INC      = 6;
parameter OP_DEC      = 7;
parameter OP_CMP      = 8;
parameter OP_ASL      = 9;
parameter OP_LSR      = 10;
parameter OP_ROL      = 11;
parameter OP_ROR      = 12;
parameter OP_UPDATE_C = 13;