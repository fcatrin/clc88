parameter OP_NOP      = 4'd0;
parameter OP_UPDATE   = 4'd1;
parameter OP_AND      = 4'd2;
parameter OP_OR       = 4'd3;
parameter OP_EOR      = 4'd4;
parameter OP_ADC      = 4'd5;
parameter OP_INC      = 4'd6;
parameter OP_DEC      = 4'd7;
parameter OP_CMP      = 4'd8;
parameter OP_ASL      = 4'd9;
parameter OP_LSR      = 4'd10;
parameter OP_ROL      = 4'd11;
parameter OP_ROR      = 4'd12;
parameter OP_BIT      = 4'd13;
parameter OP_UPDATE_C = 4'd14;